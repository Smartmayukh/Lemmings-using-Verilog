module counter (

    input clk,

    input reset,

    input areset,

    output signal);

    reg [5:0] count;
  
  

    always@(posedge clk)begin
      

        if(areset || (reset && count<6'd19) )

            begin

            count=6'd0;

            signal=0;

            end

        else if(~reset && count<6'd19)

            begin

            count++;

            signal=0;

            end

        else if(reset && count>=6'd19)

            begin

            count=6'd0;

            signal=1;

            end

        else

            signal=1;

            

    end

endmodule





module top_module(

    input clk,

    input areset,    

    input bump_left,

    input bump_right,

    input ground,

    input dig,

    output walk_left,

    output walk_right,

    output aaah,

    output digging ); 

    

    parameter LEFT=0,RIGHT=1,FALLING_LEFT=2,FALLING_RIGHT=3,DIGGING_LEFT=4,DIGGING_RIGHT=5,SPLAT=6;

    

    reg [2:0] state, next_state;

    

    wire splat_left,splat_right;

    

    counter A(clk,~(state==FALLING_LEFT),areset,splat_left);

    counter B(clk,~(state==FALLING_RIGHT),areset,splat_right);



    

    always @(*) begin

        case(state)

            LEFT:           next_state=(~ground)   ?    FALLING_LEFT   : ((dig)?  DIGGING_LEFT:((bump_left)?RIGHT:LEFT));

            RIGHT:          next_state=(~ground)   ?    FALLING_RIGHT  : ((dig)?  DIGGING_RIGHT:((bump_right )?LEFT:RIGHT));  

            FALLING_LEFT:   next_state=(ground)    ?    ((splat_left==1)? SPLAT:LEFT)  : FALLING_LEFT;

            FALLING_RIGHT:  next_state=(ground)    ?    ((splat_right==1)? SPLAT:RIGHT): FALLING_RIGHT;

            DIGGING_LEFT:   next_state=(ground)    ?    DIGGING_LEFT   : FALLING_LEFT;

            DIGGING_RIGHT:  next_state=(ground)    ?    DIGGING_RIGHT  : FALLING_RIGHT;

            SPLAT :         next_state=SPLAT;

        endcase

    end

  
  


    always @(posedge clk, posedge areset) begin

        if(areset==1)

            state<=LEFT;

        else

            state<=next_state;

    end

            

            

    assign walk_left=(state==LEFT)&&~(state==SPLAT);
  

    assign walk_right=(state==RIGHT)&&~(state==SPLAT);
  

    assign aaah=(state==FALLING_LEFT || state==FALLING_RIGHT)&&~(state==SPLAT);
  

    assign digging=(state==DIGGING_LEFT || state==DIGGING_RIGHT)&&~(state==SPLAT);           




endmodule
